library verilog;
use verilog.vl_types.all;
entity EXP_tb is
end EXP_tb;
