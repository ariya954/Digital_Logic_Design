library verilog;
use verilog.vl_types.all;
entity tb_ASSUME_R4 is
end tb_ASSUME_R4;
