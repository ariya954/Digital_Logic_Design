library verilog;
use verilog.vl_types.all;
entity Function_Generator_TestBench is
end Function_Generator_TestBench;
