library verilog;
use verilog.vl_types.all;
entity counter_Testbench is
end counter_Testbench;
