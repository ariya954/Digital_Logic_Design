`timescale 1ns/1ns

module Register(input clk, reset, load, input [19 : 0] D, output reg [19 : 0]Q);

always @(posedge clk, posedge reset)begin
   if(reset)
      Q <= 20'b0;
   else begin
      if(load)
         Q <= D;
   end
end

endmodule

module eight_bit_Decoder(input [7 : 0]_input, output reg[149 : 0]decoded_output);

reg [7 : 0]i, j;
always @(_input)begin
  for(i = 0; i < 150; i = i + 1)begin
    decoded_output[i] = 1'b0;
  end
  decoded_output[_input] = 1'b1;
end

endmodule

module Error_Checker_DataPath(input clk, reset, input [19 : 0]x_Bus, y_Bus, b_0, b_1, input [7 : 0]output_select, register_load_select, output [19 : 0]error);

wire [19 : 0] x [149 : 0];
wire [19 : 0] y [149 : 0];
wire [149 : 0]load;

eight_bit_Decoder Decoder(register_load_select, load);
genvar k;
generate
for(k = 0; k < 150; k = k + 1) 
 begin
   Register xx(clk, reset, load[k], x_Bus, x[k]); 
   Register yy(clk, reset, load[k], y_Bus, y[k]); 
 end 
endgenerate

assign error =  y[output_select] - (b_1 * x[output_select]) - b_0;

endmodule

module Error_Checker_CU(input en, clk, reset, output reg[7 : 0]register_load_select, output_select);

wire co_of_counter_of_Decoder_input, co_of_counter_of_Mux_select;
reg[2 : 0] ns, ps;
parameter[2 : 0] Idle = 3'b000, load_data = 3'b001, Inc_load = 3'b010, calculate_error = 3'b011, send_calculated_error = 3'b100;
always @(en, ps, co_of_counter_of_Decoder_input, co_of_counter_of_Mux_select) begin
   case(ps) 
     Idle:  begin ns = en ? load_data : Idle; end
     load_data:  begin ns = Inc_load; register_load_select = register_load_select + 1; end
     Inc_load: begin ns = co_of_counter_of_Decoder_input ? calculate_error : load_data; register_load_select = register_load_select + 1; end
     calculate_error: begin ns = send_calculated_error; output_select = output_select + 1; end
     send_calculated_error: begin ns = co_of_counter_of_Mux_select ? Idle : calculate_error; output_select = output_select + 1; end
     default: begin ns = Idle; register_load_select = 8'b0; output_select = 8'b0; end
   endcase
end

always @(posedge clk, posedge reset) begin
   if(reset)
     ps <= 0;
   else begin
     ps <= ns;
   end
end

assign co_of_counter_of_Decoder_input = (register_load_select >= 150) ? 1 : 0;
assign co_of_counter_of_Mux_select = (output_select >= 150) ? 1 : 0;
assign output_select = output_select < 150 ? output_select : 0;

endmodule

module Error_Checker(input en, clk, reset, input [19 : 0]b_0, b_1, x_Bus, y_Bus, output [19 : 0]error);

wire [7 : 0]register_load_select, output_select;
Error_Checker_DataPath Data_Path(clk, reset, x_Bus, y_Bus, b_0, b_1, output_select, register_load_select, error);
Error_Checker_CU CU(en, clk, reset, register_load_select, output_select);

endmodule
